module day_01

fn part_one(input string) int {
	return input.len
}
