module day_01

import os

fn test_part_one() ! {
	assert part_one(input: "Hello, World!")! == 13
}

fn test_part_two() {
	assert part_two()! == 28
}
